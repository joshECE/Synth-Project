module top_module (

);

